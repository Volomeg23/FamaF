./SingleCycleProcessor/alu.sv