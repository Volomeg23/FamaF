./SingleCycleProcessor/signext.sv