module imem #(parameter N = 32) ( // Los warnings están bien
		input logic [5:0] addr,
		output logic [N-1:0] q
	);

	logic [N-1:0] rom [0:63] = '{default: 32'h0};

	initial begin
				rom[0:127] = 
	'{32'h8b050083, 32'hf8018003, 32'hcb050083, 32'hf8020003, 32'hcb0a03e4, 32'hf8028004, 32'h8b040064, 32'hf8030004, 	
	  32'hcb030025, 32'hf8038005, 32'h8a1f0145, 32'hf8040005, 32'h8a030145, 32'hf8048005, 32'h8a140294, 32'hf8050014, 	
	  32'haa1f0166, 32'hffffffff, 32'hf8058006, 32'hf846000c, 32'hf806800c, 32'h8b1c039c, 32'h8b18039c, 32'h8b18039c, 	
	  32'h8b18039c, 32'hd61f0380, 32'hf8000001, 32'hf8008002, 32'hf8000203, 32'h00000000, 32'h00000000, 32'h00000000, 	
	  32'h8b1f03ed, 32'h8b0101ad, 32'hf807000d, 32'hb4ffffdf, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hd5382014, 32'hcb020294, 
	  32'hb4000094, 32'h8b0103bd, 32'hf808801d, 32'hd69f03e0, 32'h8b0103de, 32'hf809001e, 32'hd5380015, 32'hd61f02a0,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
	  32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
	end

	always_comb begin
		q = rom[addr];
	end

endmodule