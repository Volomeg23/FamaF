./SingleCycleProcessor/imem.sv