./SingleCycleProcessor/regfile.sv