./SingleCycleProcessor/execute.sv