./SingleCycleProcessor/maindec.sv