./SingleCycleProcessor/adder.sv