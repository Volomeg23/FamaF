./SingleCycleProcessor/mux2.sv