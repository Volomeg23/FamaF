./SingleCycleProcessor/fetch.sv