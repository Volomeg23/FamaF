./SingleCycleProcessor/flopr.sv