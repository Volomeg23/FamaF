./SingleCycleProcessor/sl2.sv